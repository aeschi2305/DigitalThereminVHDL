-- Audio.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Audio is
	port (
		to_dac_left_channel_data     : in  std_logic_vector(31 downto 0) := (others => '0'); --    avalon_left_channel_sink.data
		to_dac_left_channel_valid    : in  std_logic                     := '0';             --                            .valid
		to_dac_left_channel_ready    : out std_logic;                                        --                            .ready
		--from_adc_left_channel_ready  : in  std_logic                     := '0';             --  avalon_left_channel_source.ready
		--from_adc_left_channel_data   : out std_logic_vector(31 downto 0);                    --                            .data
		--from_adc_left_channel_valid  : out std_logic;                                        --                            .valid
		to_dac_right_channel_data    : in  std_logic_vector(31 downto 0) := (others => '0'); --   avalon_right_channel_sink.data
		to_dac_right_channel_valid   : in  std_logic                     := '0';             --                            .valid
		to_dac_right_channel_ready   : out std_logic;                                        --                            .ready
		--from_adc_right_channel_ready : in  std_logic                     := '0';             -- avalon_right_channel_source.ready
		--from_adc_right_channel_data  : out std_logic_vector(31 downto 0);                    --                            .data
		--from_adc_right_channel_valid : out std_logic;                                        --                            .valid
		clk                          : in  std_logic                     := '0';             --                         clk.clk
		AUD_BCLK                     : in  std_logic                     := '0';             --          external_interface.BCLK
		AUD_DACDAT                   : out std_logic;                                        --                            .DACDAT
		AUD_DACLRCK                  : in  std_logic                     := '0';             --                            .DACLRCK
		reset                        : in  std_logic                     := '0'              --                       reset.reset
	);
end entity Audio;

architecture rtl of Audio is
	component Audio_audio_0 is
		port (
			clk                          : in  std_logic                     := 'X';             -- clk
			reset                        : in  std_logic                     := 'X';             -- reset
			--from_adc_left_channel_ready  : in  std_logic                     := 'X';             -- ready
			--from_adc_left_channel_data   : out std_logic_vector(31 downto 0);                    -- data
			--from_adc_left_channel_valid  : out std_logic;                                        -- valid
			--from_adc_right_channel_ready : in  std_logic                     := 'X';             -- ready
			--from_adc_right_channel_data  : out std_logic_vector(31 downto 0);                    -- data
			--from_adc_right_channel_valid : out std_logic;                                        -- valid
			to_dac_left_channel_data     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			to_dac_left_channel_valid    : in  std_logic                     := 'X';             -- valid
			to_dac_left_channel_ready    : out std_logic;                                        -- ready
			to_dac_right_channel_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			to_dac_right_channel_valid   : in  std_logic                     := 'X';             -- valid
			to_dac_right_channel_ready   : out std_logic;                                        -- ready
			AUD_BCLK                     : in  std_logic                     := 'X';             -- export
			AUD_DACDAT                   : out std_logic;                                        -- export
			AUD_DACLRCK                  : in  std_logic                     := 'X'              -- export
		);
	end component Audio_audio_0;

begin

	audio_0 : component Audio_audio_0
		port map (
			clk                          => clk,                          --                         clk.clk
			reset                        => reset,                        --                       reset.reset
			--from_adc_left_channel_ready  => from_adc_left_channel_ready,  --  avalon_left_channel_source.ready
			--from_adc_left_channel_data   => from_adc_left_channel_data,   --                            .data
			--from_adc_left_channel_valid  => from_adc_left_channel_valid,  --                            .valid
			--from_adc_right_channel_ready => from_adc_right_channel_ready, -- avalon_right_channel_source.ready
			--from_adc_right_channel_data  => from_adc_right_channel_data,  --                            .data
			--from_adc_right_channel_valid => from_adc_right_channel_valid, --                            .valid
			to_dac_left_channel_data     => to_dac_left_channel_data,     --    avalon_left_channel_sink.data
			to_dac_left_channel_valid    => to_dac_left_channel_valid,    --                            .valid
			to_dac_left_channel_ready    => to_dac_left_channel_ready,    --                            .ready
			to_dac_right_channel_data    => to_dac_right_channel_data,    --   avalon_right_channel_sink.data
			to_dac_right_channel_valid   => to_dac_right_channel_valid,   --                            .valid
			to_dac_right_channel_ready   => to_dac_right_channel_ready,   --                            .ready
			AUD_BCLK                     => AUD_BCLK,                     --          external_interface.export
			AUD_DACDAT                   => AUD_DACDAT,                   --                            .export
			AUD_DACLRCK                  => AUD_DACLRCK                   --                            .export
		);

end architecture rtl; -- of Audio
