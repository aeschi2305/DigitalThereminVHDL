-- Audio_clock.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Audio_clock is
	port (
		audio_clk_clk      : out std_logic;        --    audio_clk.clk
		ref_clk_clk        : in  std_logic := '0'; --      ref_clk.clk
		ref_reset_reset    : in  std_logic := '0'; --    ref_reset.reset
		reset_source_reset : out std_logic         -- reset_source.reset
	);
end entity Audio_clock;

architecture rtl of Audio_clock is
	component Audio_clock_audio_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			audio_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component Audio_clock_audio_pll_0;

begin

	audio_pll_0 : component Audio_clock_audio_pll_0
		port map (
			ref_clk_clk        => ref_clk_clk,        --      ref_clk.clk
			ref_reset_reset    => ref_reset_reset,    --    ref_reset.reset
			audio_clk_clk      => audio_clk_clk,      --    audio_clk.clk
			reset_source_reset => reset_source_reset  -- reset_source.reset
		);

end architecture rtl; -- of Audio_clock
